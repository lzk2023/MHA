`timescale 1ns/1ps
module tb_SA_wrapper(

);
localparam D_W = 16;
localparam S   = 16;
localparam C   = 16;

bit                     I_CLK        ;
bit                     I_RST_N      ;
bit                     I_START_FLAG ;
bit                     I_END_FLAG   ;
bit   [(S*D_W)-1:0]     I_X          ;
bit   [(C*D_W)-1:0]     I_W          ;
  
logic                   O_OUT_VLD    ;
logic  [(S*C*D_W)-1:0]  O_OUT        ;
logic                   O_PE_SHIFT   ;

bit [D_W-1:0] X_MATRIX [0:S-1][0:C-1];
bit [D_W-1:0] W_MATRIX [0:S-1][0:C-1];
bit [D_W-1:0] O_MATRIX [0:S-1][0:C-1];
bit [15:0] sel;

SA_wrapper#(
    .D_W     (D_W          ),
    .S       (S            ),  //SA_ROW,        SA.shape = (S,C)
    .C       (C            )   //SA_COLUMN,     
) u_dut_SA_top(
    .I_CLK       (I_CLK        ),
    .I_RST_N     (I_RST_N      ),
    .I_START_FLAG(I_START_FLAG ),//
    .I_END_FLAG  (   ),                                                
    .I_X         (I_X          ),//input x(from left)     
    .I_W         (I_W          ),//input weight(from ddr)             
    .O_OUT_VLD   (O_OUT_VLD    ),// 
    .O_PE_SHIFT  (O_PE_SHIFT   ),                                  
    .O_OUT       (O_OUT        ) //OUT.shape = (X_R,64)               
);           

always #5 I_CLK = ~I_CLK;
generate 
    for(genvar i=0;i<S;i=i+1)begin
        assign I_X[i*D_W +: D_W] = X_MATRIX[i][S-1-sel];
    end
endgenerate

generate 
    for(genvar i=0;i<C;i=i+1)begin
        assign I_W[i*D_W +: D_W] = W_MATRIX[S-1-sel][i];
    end
endgenerate

generate 
    for(genvar i=0;i<S;i=i+1)begin
        for(genvar j=0;j<C;j=j+1)begin
            assign O_MATRIX[i][j] = O_OUT[(i*C+j)*D_W +: D_W];
        end
    end
endgenerate
always@(posedge I_CLK or negedge I_RST_N)begin
    if(!I_RST_N)begin
        sel <= 0;
    end else if(O_PE_SHIFT)begin
        if(sel<S-1)begin
            sel <= sel + 1;
        end else begin
            sel <= sel;
        end
    end
end

//function [15:0] mul_16;
//    input [15:0] a;
//    input [15:0] b;
//    reg [31:0] c;
//    begin
//        c = $signed(a) * $signed(b);
//        mul_16 = {c[31],c[27:13]};
//    end
//endfunction

initial begin
    #100
    I_RST_N = 1;
    I_START_FLAG = 1;
    X_MATRIX = '{
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00}
    };
    W_MATRIX = '{
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00},
        '{16'h000,16'h100,16'h200,16'h300,16'h400,16'h500,16'h600,16'h700,16'h800,16'h900,16'ha00,16'hb00,16'hc00,16'hd00,16'he00,16'hf00}
    };
    //X_MATRIX = '{
    //    '{16'h000,16'h100,16'h200},
    //    '{16'h000,16'h100,16'h200},
    //    '{16'h000,16'h100,16'h200}
    //};
    //W_MATRIX = '{
    //    '{16'h000,16'h100,16'h200},
    //    '{16'h000,16'h100,16'h200},
    //    '{16'h000,16'h100,16'h200}
    //};
    #10
    I_START_FLAG = 0;
    #50000
    $finish;
end
endmodule
