`timescale 1ns/1ps
module flash_attn();
endmodule