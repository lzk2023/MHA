`timescale 1ns/1ps
module flash_attn_top(
    input  logic        I_CLK  ,
    input  logic        I_RST_N,
    input  logic        I_START,
    output logic        O_VLD  ,
    output logic [15:0] O_OUT  
);

endmodule