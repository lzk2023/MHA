`timescale 1ns/1ps
module bram_mi_li(
    input  logic       I_CLK             , 
    input  logic       I_RST_N           , 
    input  logic       I_RD_ENA          ,
    input  logic       I_WR_ENA          
);

endmodule